--
-- VHDL Architecture ece411.Memory.UNTITLED
--
-- Created:
--          by - baker30.ews (siebl-0220-06.ews.illinois.edu)
--          at - 04:22:04 01/22/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Memory IS
   PORT( 
      ADDRESS   : IN     LC3b_word;
      DATAOUT   : IN     LC3b_word;
      MREAD_L   : IN     std_logic;
      MWRITEH_L : IN     std_logic;
      MWRITEL_L : IN     std_logic;
      RESET_L   : IN     std_logic;
      clk       : IN     std_logic;
      DATAIN    : OUT    LC3b_word;
      MRESP_H   : OUT    std_logic
   );

-- Declarations

END Memory ;

--
-- VHDL Architecture ece411.Memory.struct
--
-- Created:
--          by - baker30.ews (evrt-252-27.ews.illinois.edu)
--          at - 17:49:11 03/03/13
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;


ARCHITECTURE struct OF Memory IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL CacheWrite : std_logic;
   SIGNAL DirtyOut   : std_logic;
   SIGNAL Evict_H    : std_logic;
   SIGNAL LRUOut     : std_logic;
   SIGNAL PMADDRESS  : LC3B_WORD;
   SIGNAL PMDATAIN   : LC3B_OWORD;
   SIGNAL PMDATAOUT  : LC3B_OWORD;
   SIGNAL PMREAD_L   : STD_LOGIC;
   SIGNAL PMRESP_H   : STD_LOGIC;
   SIGNAL PMWRITE_L  : STD_LOGIC;
   SIGNAL hit        : std_logic;


   -- Component Declarations
   COMPONENT Cache_Controller
   PORT (
      DirtyOut   : IN     std_logic ;
      LRUOut     : IN     std_logic ;
      MWRITEL_L  : IN     std_logic ;
      PMRESP_H   : IN     STD_LOGIC ;
      RESET_L    : IN     std_logic ;
      clk        : IN     std_logic ;
      hit        : IN     std_logic ;
      CacheWrite : OUT    std_logic ;
      Evict_H    : OUT    std_logic ;
      PMREAD_L   : OUT    STD_LOGIC ;
      PMWRITE_L  : OUT    STD_LOGIC 
   );
   END COMPONENT;
   COMPONENT Cache_Datapath
   PORT (
      ADDRESS    : IN     LC3b_word ;
      CacheWrite : IN     std_logic ;
      DATAOUT    : IN     LC3b_word ;
      Evict_H    : IN     std_logic ;
      MREAD_L    : IN     std_logic ;
      MWRITEH_L  : IN     std_logic ;
      MWRITEL_L  : IN     std_logic ;
      PMDATAIN   : IN     LC3B_OWORD ;
      RESET_L    : IN     std_logic ;
      clk        : IN     std_logic ;
      DATAIN     : OUT    LC3b_word ;
      DirtyOut   : OUT    std_logic ;
      LRUOut     : OUT    std_logic ;
      MRESP_H    : OUT    std_logic ;
      PMADDRESS  : OUT    LC3B_WORD ;
      PMDATAOUT  : OUT    LC3B_OWORD ;
      hit        : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Physical_Memory
   PORT (
      clk       : IN     std_logic ;
      PMADDRESS : IN     LC3B_WORD ;
      PMDATAOUT : IN     LC3B_OWORD ;
      PMREAD_L  : IN     STD_LOGIC ;
      RESET_L   : IN     std_logic ;
      PMDATAIN  : OUT    LC3B_OWORD ;
      PMRESP_H  : OUT    STD_LOGIC ;
      PMWRITE_L : IN     STD_LOGIC 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Cache_Controller USE ENTITY ece411.Cache_Controller;
   FOR ALL : Cache_Datapath USE ENTITY ece411.Cache_Datapath;
   FOR ALL : Physical_Memory USE ENTITY ece411.Physical_Memory;
   -- pragma synthesis_on


BEGIN

   -- Instance port mappings.
   Cache_Cont : Cache_Controller
      PORT MAP (
         DirtyOut   => DirtyOut,
         LRUOut     => LRUOut,
         MWRITEL_L  => MWRITEL_L,
         PMRESP_H   => PMRESP_H,
         RESET_L    => RESET_L,
         clk        => clk,
         hit        => hit,
         CacheWrite => CacheWrite,
         Evict_H    => Evict_H,
         PMREAD_L   => PMREAD_L,
         PMWRITE_L  => PMWRITE_L
      );
   Cache_DP : Cache_Datapath
      PORT MAP (
         ADDRESS    => ADDRESS,
         CacheWrite => CacheWrite,
         DATAOUT    => DATAOUT,
         Evict_H    => Evict_H,
         MREAD_L    => MREAD_L,
         MWRITEH_L  => MWRITEH_L,
         MWRITEL_L  => MWRITEL_L,
         PMDATAIN   => PMDATAIN,
         RESET_L    => RESET_L,
         clk        => clk,
         DATAIN     => DATAIN,
         DirtyOut   => DirtyOut,
         LRUOut     => LRUOut,
         MRESP_H    => MRESP_H,
         PMADDRESS  => PMADDRESS,
         PMDATAOUT  => PMDATAOUT,
         hit        => hit
      );
   PDRAM : Physical_Memory
      PORT MAP (
         clk       => clk,
         PMADDRESS => PMADDRESS,
         PMDATAOUT => PMDATAOUT,
         PMREAD_L  => PMREAD_L,
         RESET_L   => RESET_L,
         PMDATAIN  => PMDATAIN,
         PMRESP_H  => PMRESP_H,
         PMWRITE_L => PMWRITE_L
      );

END struct;
